`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    10:32:26 11/07/2016 
// Design Name: 
// Module Name:    MemoriaParaIntrucciones 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module MemoriaParaIntrucciones(
	 input [31:0] address,
    output reg [31:0] dataOutput
    );
	 
	 always@*
	 begin                                            
		case(address)
				32'h00:      dataOutput = 32'b11100010000010011001111100000000 ; 
				/*------------Logica de espera------*/
				32'h04:      dataOutput = 32'b11100010000010011001111100000000 ;  
				32'h08:      dataOutput = 32'b11100010000000000000111100000000 ;   
				32'h0C:      dataOutput = 32'b11100010000000110011111100000000 ;  
				32'h10:      dataOutput = 32'b11100010100010011001111100010000 ;  
				32'h14:      dataOutput = 32'b11100101101110010001000000000000 ;  
				32'h18:      dataOutput = 32'b11100101101110010010000000000100 ;
				32'h1C:      dataOutput = 32'b11100101101110111101000000000000 ;     
				32'h20:      dataOutput = 32'b11100011010111011111111100000001 ;
				32'h24:      dataOutput = 32'b00001010000000000000000000001001 ;
				32'h28:      dataOutput = 32'b11100011010111011111111100000010 ;
				32'h2C:      dataOutput = 32'b00001010000000000000000000001111 ;
				32'h30:      dataOutput = 32'b11100011010111011111111100000011 ;
				32'h34:      dataOutput = 32'b00001010000000000000000000010001 ;
				32'h38:      dataOutput = 32'b11100011010111011111111100000100 ;
				32'h3C:      dataOutput = 32'b00001010000000000000000000010011 ;
				32'h40:      dataOutput = 32'b11100011010111011111111100000101 ;
				32'h44:      dataOutput = 32'b00001010000000000000000000011011 ;
				32'h48:      dataOutput = 32'b11100011010111011111111100000000 ;               
				32'h4C:      dataOutput = 32'b11101010111111111111111111101100 ;
							/*------------MULTIPLICACION------*/
				32'h50:      dataOutput = 32'b11100011100011001100111100000001 ;
				32'h54:      dataOutput = 32'b11100001010100101111000000000011 ;       
				32'h58:      dataOutput = 32'b00010000100000000000000000000001 ;         
				32'h5C:      dataOutput = 32'b00010000100000110011000000001100 ;          
				32'h60:      dataOutput = 32'b00011010111111111111111111111011 ;                                     
				32'h64:      dataOutput = 32'b11100101101010010000000000001000 ;        
				32'h68:      dataOutput = 32'b11100010000011011101111100000000 ;
				32'h6C:      dataOutput = 32'b11101010111111111111111111100100 ;  
									
									/*------------SUMA-----------*/
					
				32'h70:    	dataOutput = 32'b11100000100000010000000000000010 ;
				32'h74:    	dataOutput = 32'b11100101101010010000000000001000 ;          
				32'h78:   	dataOutput = 32'b11100010000011011101111100000000 ;
				32'h7c:     dataOutput = 32'b11101010111111111111111111100000 ;
								  
								  /*------------RESTA-----------*/
						
				32'h80:    	dataOutput = 32'b11100000010000010000000000000010 ;
				32'h84:    	dataOutput = 32'b11100101101010010000000000001000 ;          
				32'h88:   	dataOutput = 32'b11100010000011011101111100000000 ;
				32'h8c:     dataOutput = 32'b11101010111111111111111111011100 ;
						 
								 /*-----------------------------DIVISION---------------------*/
								 
									
				32'h90:      dataOutput = 32'b11100011100011001100111100000001 ;
				32'h94:      dataOutput = 32'b11100011010100101111111100000000 ; 
				32'h98:      dataOutput = 32'b00001010111111111111111111011100 ;         
				32'h9C:      dataOutput = 32'b11100001010100101111000000000001 ;           
				32'hA0:      dataOutput = 32'b10010000100000000000111111111100 ;           
				32'hA4:      dataOutput = 32'b10010000010000010001111111110010 ;         
				32'hA8:      dataOutput = 32'b10011010111111111111111111111011 ;          
				32'hAC:      dataOutput = 32'b11100101101010010000000000001000 ;    
				32'hB0: 	 dataOutput = 32'b11100010000011011101111100000000 ;
				32'hB4:      dataOutput = 32'b11101010111111111111111111010010 ;
						  
									/*-----------------------------MODULO---------------------*/
									 
				32'hB8:      dataOutput = 32'b11100011010100101111111100000000 ; 
				32'hBC:      dataOutput = 32'b00001010000000000000000000000010 ;
				32'hC0:      dataOutput = 32'b11100001010100101111111111110001 ;
				32'hC4:      dataOutput = 32'b10010000010000010001111111110010 ;
				32'hC8:      dataOutput = 32'b10011010111111111111111111111100 ;
				32'hCC:      dataOutput = 32'b11100001100000010000111111110000 ;
				32'hD0:      dataOutput = 32'b11100101101010010000000000001000 ;   
				32'hD4:      dataOutput = 32'b11100010000011011101111100000000 ;
				32'hD8:      dataOutput = 32'b11101010111111111111111111001001 ;
				
		
				default: dataOutput = 32'b0;
		endcase
	 end
endmodule
